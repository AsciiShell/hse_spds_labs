
module de0_cv
(
    input           CLOCK2_50,
    input           CLOCK3_50,
    inout           CLOCK4_50,
    input           CLOCK_50,
                   
    input           RESET_N,

    input   [ 3:0]  KEY,
    input   [ 9:0]  SW,

    output  [ 9:0]  LEDR,

    output  [ 6:0]  HEX0,
    output  [ 6:0]  HEX1,
    output  [ 6:0]  HEX2,
    output  [ 6:0]  HEX3,
    output  [ 6:0]  HEX4,
    output  [ 6:0]  HEX5,
                   
    output  [12:0]  DRAM_ADDR,
    output  [ 1:0]  DRAM_BA,
    output          DRAM_CAS_N,
    output          DRAM_CKE,
    output          DRAM_CLK,
    output          DRAM_CS_N,
    inout   [15:0]  DRAM_DQ,
    output          DRAM_LDQM,
    output          DRAM_RAS_N,
    output          DRAM_UDQM,
    output          DRAM_WE_N,
                   
    output  [ 3:0]  VGA_B,
    output  [ 3:0]  VGA_G,
    output          VGA_HS,
    output  [ 3:0]  VGA_R,
    output          VGA_VS,

    inout           PS2_CLK,
    inout           PS2_CLK2,
    inout           PS2_DAT,
    inout           PS2_DAT2,
                   
    output          SD_CLK,
    inout           SD_CMD,
    inout   [ 3:0]  SD_DATA,
                   
    inout   [35:0]  GPIO_0,
    inout   [35:0]  GPIO_1
);

    // wires & inputs
    wire          clk;
    wire          clkIn     =  CLOCK_50;
    wire          rst_n     =  KEY[0] & RESET_N;
    wire          clkEnable =  SW [9] | ~KEY[1];
    wire [  3:0 ] clkDevide =  SW [8:5];
    wire [  4:0 ] regAddr   =  SW [4:0];
    wire [ 31:0 ] regData;
    wire [ `SM_GPIO_WIDTH - 1:0] gpioInput = { 8'b0, GPIO_0 [7:0]};
	 wire [ `SM_GPIO_WIDTH - 1:0] gpioOutput;

    //cores
    sm_top sm_top
    (
        .clkIn      ( clkIn     ),
        .rst_n      ( rst_n     ),
        .clkDevide  ( clkDevide ),
        .clkEnable  ( clkEnable ),
        .clk        ( clk       ),
        .regAddr    ( regAddr   ),
        .regData    ( regData   ),
        .gpioInput  ( gpioInput ),
        .gpioOutput ( gpioOutput)
    );

    //outputs
    assign LEDR[0]   = clk;
    assign LEDR[9:1] = regData[8:0];

    wire [ 31:0 ] h7segment = regData;

    sm_hex_display digit_5 ( GPIO_0 [7:4] , HEX5 [6:0] );
    sm_hex_display digit_4 ( GPIO_0 [3:0] , HEX4 [6:0] );
    sm_hex_display digit_3 ( h7segment [15:12] , HEX3 [6:0] );
    sm_hex_display digit_2 ( h7segment [11: 8] , HEX2 [6:0] );
    sm_hex_display digit_1 ( h7segment [ 7: 4] , HEX1 [6:0] );
    sm_hex_display digit_0 ( h7segment [ 3: 0] , HEX0 [6:0] );

    wire [15:0] h7segment_my = 4'habcd;
    wire [6:0] digit1;
    wire [6:0] digit2;
    wire [6:0] digit3;
	 //wire [11:0] gpio1;
    //assign GPIO_1 [11:0] = gpio1[11:0];
    sm_hex_display_our digit_2_our ( h7segment_my [11: 8] , digit1 [6:0] );
    sm_hex_display_our digit_1_our ( h7segment_my [ 7: 4] , digit2 [6:0] );
    sm_hex_display_our digit_0_our ( h7segment_my [ 3: 0] , digit3 [6:0] );
    sm_hex_display_digit dis_digit (
        .digit1 (digit1),
        .digit2 (digit2),
        .digit3 (digit3),
        .clkIn  (clkIn),
        .seven_segments (GPIO_1 [11:0])
    );

endmodule
