module SEG7_LUT_6 (	oSEG0,oSEG1,oSEG2,oSEG3,oSEG4,oSEG5,iDIG , key);
input	[23:0]	iDIG;
input				key;
output	[6:0]	oSEG0,oSEG1,oSEG2,oSEG3,oSEG4,oSEG5;

//SEG7_LUT	u0	(	oSEG0,iDIG[3:0]		);
//SEG7_LUT	u1	(	oSEG1,iDIG[7:4]		);
//SEG7_LUT	u2	(	oSEG2,iDIG[11:8]	);
//SEG7_LUT	u3	(	oSEG3,iDIG[15:12]	);
//SEG7_LUT	u4	(	oSEG4,iDIG[19:16]	);
//SEG7_LUT	u5	(	oSEG5,iDIG[23:20]	);

SEG7_LUT_m	u0	(	oSEG0, key, iDIG[3:0]		);
SEG7_LUT_m	u1	(	oSEG1, key, iDIG[7:4]		);
SEG7_LUT_m	u2	(	oSEG2, key, iDIG[11:8]	);
SEG7_LUT_m	u3	(	oSEG3, key, iDIG[15:12]	);
SEG7_LUT_m	u4	(	oSEG4, key, iDIG[19:16]	);
SEG7_LUT_m	u5	(	oSEG5, key, iDIG[23:20]	);


endmodule